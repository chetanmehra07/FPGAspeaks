module not_1(in,out);
  input in;
  output out;
  assign out= ~in;
endmodule
